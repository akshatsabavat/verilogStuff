`timescale 1ps/1ns
`include "hello.v"

module hello_tb():
    reg A, B;
    hello_uut(A,B);

    initial begin
        $dumpfile("hello_tb.vcd")
        $dumpvars(0, hello_tb)

        A = 0;
        #20;

        A = 1;
        #20;

        A=0;
        #20;
    end
endmodule